--------------------------------------------------------------------------------
--  Module  : connections.vhdl
--  Author  : Andy
--  Created : April 17, 2007, 11:02 PM
--------------------------------------------------------------------------------

package connections is
  
   
end package connections;  



package body connections is

 
end package body;
